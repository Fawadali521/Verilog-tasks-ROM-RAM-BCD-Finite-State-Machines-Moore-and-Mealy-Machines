library verilog;
use verilog.vl_types.all;
entity mux2 is
end mux2;
