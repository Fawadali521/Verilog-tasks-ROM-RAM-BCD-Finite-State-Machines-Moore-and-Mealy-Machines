library verilog;
use verilog.vl_types.all;
entity stim9 is
end stim9;
