library verilog;
use verilog.vl_types.all;
entity light_test is
end light_test;
