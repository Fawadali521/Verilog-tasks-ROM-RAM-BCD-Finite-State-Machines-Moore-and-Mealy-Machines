library verilog;
use verilog.vl_types.all;
entity stim1 is
end stim1;
