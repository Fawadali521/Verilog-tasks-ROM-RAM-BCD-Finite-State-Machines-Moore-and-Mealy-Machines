library verilog;
use verilog.vl_types.all;
entity mux4 is
end mux4;
