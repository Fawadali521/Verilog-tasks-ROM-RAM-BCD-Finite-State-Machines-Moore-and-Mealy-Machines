library verilog;
use verilog.vl_types.all;
entity lock_test is
end lock_test;
