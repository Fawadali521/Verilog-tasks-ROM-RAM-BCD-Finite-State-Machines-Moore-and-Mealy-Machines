library verilog;
use verilog.vl_types.all;
entity pulse is
end pulse;
