library verilog;
use verilog.vl_types.all;
entity top_de is
end top_de;
