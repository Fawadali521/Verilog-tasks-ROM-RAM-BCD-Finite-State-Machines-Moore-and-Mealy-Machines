library verilog;
use verilog.vl_types.all;
entity st is
end st;
