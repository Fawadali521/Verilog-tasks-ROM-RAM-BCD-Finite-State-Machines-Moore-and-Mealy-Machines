library verilog;
use verilog.vl_types.all;
entity stim6 is
end stim6;
