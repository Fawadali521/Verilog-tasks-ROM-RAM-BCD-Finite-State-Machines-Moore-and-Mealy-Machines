module buffer(a,b); 
input a;
output b; 
buf x1(a,b); 
endmodule
