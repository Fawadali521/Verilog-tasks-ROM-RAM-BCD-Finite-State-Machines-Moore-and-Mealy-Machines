library verilog;
use verilog.vl_types.all;
entity railway_test is
end railway_test;
