library verilog;
use verilog.vl_types.all;
entity stim5 is
end stim5;
