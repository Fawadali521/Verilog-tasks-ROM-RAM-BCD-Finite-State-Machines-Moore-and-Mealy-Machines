library verilog;
use verilog.vl_types.all;
entity stim4 is
end stim4;
