library verilog;
use verilog.vl_types.all;
entity swith is
end swith;
