library verilog;
use verilog.vl_types.all;
entity mux21_test is
end mux21_test;
