library verilog;
use verilog.vl_types.all;
entity tst_parity_rst is
end tst_parity_rst;
