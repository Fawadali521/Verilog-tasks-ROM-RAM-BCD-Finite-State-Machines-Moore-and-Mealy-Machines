library verilog;
use verilog.vl_types.all;
entity tst_moore is
end tst_moore;
