library verilog;
use verilog.vl_types.all;
entity tst_mealy is
end tst_mealy;
