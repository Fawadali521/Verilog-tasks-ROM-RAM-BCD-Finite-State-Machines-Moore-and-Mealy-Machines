library verilog;
use verilog.vl_types.all;
entity stim7 is
end stim7;
