library verilog;
use verilog.vl_types.all;
entity test_led is
end test_led;
