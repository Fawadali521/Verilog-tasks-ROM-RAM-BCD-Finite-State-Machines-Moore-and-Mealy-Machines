library verilog;
use verilog.vl_types.all;
entity stim8 is
end stim8;
