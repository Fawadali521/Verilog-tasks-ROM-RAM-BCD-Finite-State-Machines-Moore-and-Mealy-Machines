library verilog;
use verilog.vl_types.all;
entity stimulusbcd is
end stimulusbcd;
